// DE0_LT24_SOPC.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module DE0_LT24_SOPC (
		input  wire        alt_pll_areset_conduit_export,               //               alt_pll_areset_conduit.export
		output wire        alt_pll_c1_clk,                              //                           alt_pll_c1.clk
		output wire        alt_pll_c3_clk,                              //                           alt_pll_c3.clk
		output wire        alt_pll_locked_conduit_export,               //               alt_pll_locked_conduit.export
		output wire        alt_pll_phasedone_conduit_export,            //            alt_pll_phasedone_conduit.export
		input  wire [12:0] background_mem_s2_address,                   //                    background_mem_s2.address
		input  wire        background_mem_s2_chipselect,                //                                     .chipselect
		input  wire        background_mem_s2_clken,                     //                                     .clken
		input  wire        background_mem_s2_write,                     //                                     .write
		output wire [15:0] background_mem_s2_readdata,                  //                                     .readdata
		input  wire [15:0] background_mem_s2_writedata,                 //                                     .writedata
		input  wire [1:0]  background_mem_s2_byteenable,                //                                     .byteenable
		input  wire        clk_clk,                                     //                                  clk.clk
		input  wire        cyclonespi_spi_interface_SPI_clk,            //             cyclonespi_spi_interface.SPI_clk
		input  wire        cyclonespi_spi_interface_SPI_CS,             //                                     .SPI_CS
		input  wire        cyclonespi_spi_interface_SPI_SDI,            //                                     .SPI_SDI
		output wire        cyclonespi_spi_interface_SPI_SDO,            //                                     .SPI_SDO
		output wire [7:0]  cyclonespi_spi_interface_data_out,           //                                     .data_out
		output wire        cyclonespi_spi_interface_data_out_enable,    //                                     .data_out_enable
		output wire [7:0]  cyclonespi_spi_interface_config,             //                                     .config
		output wire        cyclonespi_spi_interface_spi_irq,            //                                     .spi_irq
		input  wire        from_key_export,                             //                             from_key.export
		input  wire        gsensor_int_external_connection_export,      //      gsensor_int_external_connection.export
		inout  wire        gsensor_spi_conduit_end_SDIO,                //              gsensor_spi_conduit_end.SDIO
		output wire        gsensor_spi_conduit_end_SCLK,                //                                     .SCLK
		output wire        gsensor_spi_conduit_end_CS_n,                //                                     .CS_n
		output wire        lt24_buffer_flag_external_connection_export, // lt24_buffer_flag_external_connection.export
		output wire        lt24_conduit_cs,                             //                         lt24_conduit.cs
		output wire        lt24_conduit_rs,                             //                                     .rs
		output wire        lt24_conduit_rd,                             //                                     .rd
		output wire        lt24_conduit_wr,                             //                                     .wr
		output wire [15:0] lt24_conduit_data,                           //                                     .data
		input  wire        lt24_conduit_0_finish_flag,                  //                       lt24_conduit_0.finish_flag
		input  wire [31:0] lt24_conduit_0_counter,                      //                                     .counter
		output wire [11:0] lt24_conduit_0_pattern,                      //                                     .pattern
		output wire [31:0] lt24_conduit_0_vx,                           //                                     .vx
		output wire [31:0] lt24_conduit_0_vy,                           //                                     .vy
		output wire [31:0] lt24_conduit_0_lt24_coin_x0,                 //                                     .lt24_coin_x0
		output wire [31:0] lt24_conduit_0_lt42_coin_y0,                 //                                     .lt42_coin_y0
		input  wire [31:0] lt24_conduit_0_lt24_coinx,                   //                                     .lt24_coinx
		input  wire [31:0] lt24_conduit_0_lt24_coin_y,                  //                                     .lt24_coin_y
		output wire [31:0] lt24_conduit_0_lt24_coin_vx0,                //                                     .lt24_coin_vx0
		output wire [31:0] lt24_conduit_0_lt24_coin_vy0,                //                                     .lt24_coin_vy0
		output wire        lt24_lcd_rstn_export,                        //                        lt24_lcd_rstn.export
		input  wire        lt24_touch_busy_export,                      //                      lt24_touch_busy.export
		input  wire        lt24_touch_penirq_n_export,                  //                  lt24_touch_penirq_n.export
		input  wire        lt24_touch_spi_MISO,                         //                       lt24_touch_spi.MISO
		output wire        lt24_touch_spi_MOSI,                         //                                     .MOSI
		output wire        lt24_touch_spi_SCLK,                         //                                     .SCLK
		output wire        lt24_touch_spi_SS_n,                         //                                     .SS_n
		input  wire [12:0] pic_mem_s2_address,                          //                           pic_mem_s2.address
		input  wire        pic_mem_s2_chipselect,                       //                                     .chipselect
		input  wire        pic_mem_s2_clken,                            //                                     .clken
		input  wire        pic_mem_s2_write,                            //                                     .write
		output wire [15:0] pic_mem_s2_readdata,                         //                                     .readdata
		input  wire [15:0] pic_mem_s2_writedata,                        //                                     .writedata
		input  wire [1:0]  pic_mem_s2_byteenable,                       //                                     .byteenable
		input  wire        reset_reset_n,                               //                                reset.reset_n
		output wire [12:0] sdram_controler_wire_addr,                   //                 sdram_controler_wire.addr
		output wire [1:0]  sdram_controler_wire_ba,                     //                                     .ba
		output wire        sdram_controler_wire_cas_n,                  //                                     .cas_n
		output wire        sdram_controler_wire_cke,                    //                                     .cke
		output wire        sdram_controler_wire_cs_n,                   //                                     .cs_n
		inout  wire [15:0] sdram_controler_wire_dq,                     //                                     .dq
		output wire [1:0]  sdram_controler_wire_dqm,                    //                                     .dqm
		output wire        sdram_controler_wire_ras_n,                  //                                     .ras_n
		output wire        sdram_controler_wire_we_n,                   //                                     .we_n
		output wire [7:0]  to_led_export                                //                               to_led.export
	);

	wire         alt_pll_c0_clk;                                               // ALT_PLL:c0 -> [CPU:clk, JTAG_UART:clk, LT24_CTRL:clk, LT24_LCD_RSTN:clk, LT24_TOUCH_BUSY:clk, LT24_TOUCH_PENIRQ_N:clk, LT24_TOUCH_SPI:clk, SDRAM_Controler:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, irq_synchronizer_004:sender_clk, mm_interconnect_0:ALT_PLL_c0_clk, rst_controller_001:clk]
	wire         alt_pll_c2_clk;                                               // ALT_PLL:c2 -> [KEY:clk, LED_CTRL:CLK, TIMER:clk, irq_synchronizer_002:receiver_clk, mm_interconnect_0:ALT_PLL_c2_clk, rst_controller_002:clk]
	wire  [31:0] cpu_data_master_readdata;                                     // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                                  // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                                  // CPU:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [26:0] cpu_data_master_address;                                      // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                   // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                         // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_readdatavalid;                                // mm_interconnect_0:CPU_data_master_readdatavalid -> CPU:d_readdatavalid
	wire         cpu_data_master_write;                                        // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                    // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                              // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                           // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                               // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                                  // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                         // mm_interconnect_0:CPU_instruction_master_readdatavalid -> CPU:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;     // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;       // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;    // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;        // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;           // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;          // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;      // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire         mm_interconnect_0_lt24_ctrl_avalon_slave_0_chipselect;        // mm_interconnect_0:LT24_CTRL_avalon_slave_0_chipselect -> LT24_CTRL:s_chipselect_n
	wire   [0:0] mm_interconnect_0_lt24_ctrl_avalon_slave_0_address;           // mm_interconnect_0:LT24_CTRL_avalon_slave_0_address -> LT24_CTRL:s_address
	wire         mm_interconnect_0_lt24_ctrl_avalon_slave_0_write;             // mm_interconnect_0:LT24_CTRL_avalon_slave_0_write -> LT24_CTRL:s_write_n
	wire  [31:0] mm_interconnect_0_lt24_ctrl_avalon_slave_0_writedata;         // mm_interconnect_0:LT24_CTRL_avalon_slave_0_writedata -> LT24_CTRL:s_writedata
	wire  [31:0] mm_interconnect_0_led_ctrl_avalon_slave_0_readdata;           // LED_CTRL:RDATA -> mm_interconnect_0:LED_CTRL_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_led_ctrl_avalon_slave_0_address;            // mm_interconnect_0:LED_CTRL_avalon_slave_0_address -> LED_CTRL:ADDR
	wire         mm_interconnect_0_led_ctrl_avalon_slave_0_read;               // mm_interconnect_0:LED_CTRL_avalon_slave_0_read -> LED_CTRL:READ
	wire         mm_interconnect_0_led_ctrl_avalon_slave_0_write;              // mm_interconnect_0:LED_CTRL_avalon_slave_0_write -> LED_CTRL:WRITE
	wire  [31:0] mm_interconnect_0_led_ctrl_avalon_slave_0_writedata;          // mm_interconnect_0:LED_CTRL_avalon_slave_0_writedata -> LED_CTRL:WDATA
	wire  [31:0] mm_interconnect_0_cyclonespi_avs_s0_readdata;                 // cycloneSPI:avs_s0_readdata -> mm_interconnect_0:cycloneSPI_avs_s0_readdata
	wire         mm_interconnect_0_cyclonespi_avs_s0_waitrequest;              // cycloneSPI:avs_s0_waitrequest -> mm_interconnect_0:cycloneSPI_avs_s0_waitrequest
	wire   [7:0] mm_interconnect_0_cyclonespi_avs_s0_address;                  // mm_interconnect_0:cycloneSPI_avs_s0_address -> cycloneSPI:avs_s0_address
	wire         mm_interconnect_0_cyclonespi_avs_s0_read;                     // mm_interconnect_0:cycloneSPI_avs_s0_read -> cycloneSPI:avs_s0_read
	wire         mm_interconnect_0_cyclonespi_avs_s0_write;                    // mm_interconnect_0:cycloneSPI_avs_s0_write -> cycloneSPI:avs_s0_write
	wire  [31:0] mm_interconnect_0_cyclonespi_avs_s0_writedata;                // mm_interconnect_0:cycloneSPI_avs_s0_writedata -> cycloneSPI:avs_s0_writedata
	wire  [31:0] mm_interconnect_0_lt24_interface_irq_0_avs_s0_readdata;       // LT24_interface_irq_0:avs_s0_readdata -> mm_interconnect_0:LT24_interface_irq_0_avs_s0_readdata
	wire         mm_interconnect_0_lt24_interface_irq_0_avs_s0_waitrequest;    // LT24_interface_irq_0:avs_s0_waitrequest -> mm_interconnect_0:LT24_interface_irq_0_avs_s0_waitrequest
	wire   [7:0] mm_interconnect_0_lt24_interface_irq_0_avs_s0_address;        // mm_interconnect_0:LT24_interface_irq_0_avs_s0_address -> LT24_interface_irq_0:avs_s0_address
	wire         mm_interconnect_0_lt24_interface_irq_0_avs_s0_read;           // mm_interconnect_0:LT24_interface_irq_0_avs_s0_read -> LT24_interface_irq_0:avs_s0_read
	wire         mm_interconnect_0_lt24_interface_irq_0_avs_s0_write;          // mm_interconnect_0:LT24_interface_irq_0_avs_s0_write -> LT24_interface_irq_0:avs_s0_write
	wire  [31:0] mm_interconnect_0_lt24_interface_irq_0_avs_s0_writedata;      // mm_interconnect_0:LT24_interface_irq_0_avs_s0_writedata -> LT24_interface_irq_0:avs_s0_writedata
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;             // CPU:jtag_debug_module_readdata -> mm_interconnect_0:CPU_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;          // CPU:jtag_debug_module_waitrequest -> mm_interconnect_0:CPU_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;          // mm_interconnect_0:CPU_jtag_debug_module_debugaccess -> CPU:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;              // mm_interconnect_0:CPU_jtag_debug_module_address -> CPU:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                 // mm_interconnect_0:CPU_jtag_debug_module_read -> CPU:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;           // mm_interconnect_0:CPU_jtag_debug_module_byteenable -> CPU:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                // mm_interconnect_0:CPU_jtag_debug_module_write -> CPU:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;            // mm_interconnect_0:CPU_jtag_debug_module_writedata -> CPU:jtag_debug_module_writedata
	wire  [31:0] mm_interconnect_0_alt_pll_pll_slave_readdata;                 // ALT_PLL:readdata -> mm_interconnect_0:ALT_PLL_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_alt_pll_pll_slave_address;                  // mm_interconnect_0:ALT_PLL_pll_slave_address -> ALT_PLL:address
	wire         mm_interconnect_0_alt_pll_pll_slave_read;                     // mm_interconnect_0:ALT_PLL_pll_slave_read -> ALT_PLL:read
	wire         mm_interconnect_0_alt_pll_pll_slave_write;                    // mm_interconnect_0:ALT_PLL_pll_slave_write -> ALT_PLL:write
	wire  [31:0] mm_interconnect_0_alt_pll_pll_slave_writedata;                // mm_interconnect_0:ALT_PLL_pll_slave_writedata -> ALT_PLL:writedata
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                            // KEY:readdata -> mm_interconnect_0:KEY_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                             // mm_interconnect_0:KEY_s1_address -> KEY:address
	wire         mm_interconnect_0_timer_s1_chipselect;                        // mm_interconnect_0:TIMER_s1_chipselect -> TIMER:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                          // TIMER:readdata -> mm_interconnect_0:TIMER_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                           // mm_interconnect_0:TIMER_s1_address -> TIMER:address
	wire         mm_interconnect_0_timer_s1_write;                             // mm_interconnect_0:TIMER_s1_write -> TIMER:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                         // mm_interconnect_0:TIMER_s1_writedata -> TIMER:writedata
	wire         mm_interconnect_0_lt24_lcd_rstn_s1_chipselect;                // mm_interconnect_0:LT24_LCD_RSTN_s1_chipselect -> LT24_LCD_RSTN:chipselect
	wire  [31:0] mm_interconnect_0_lt24_lcd_rstn_s1_readdata;                  // LT24_LCD_RSTN:readdata -> mm_interconnect_0:LT24_LCD_RSTN_s1_readdata
	wire   [1:0] mm_interconnect_0_lt24_lcd_rstn_s1_address;                   // mm_interconnect_0:LT24_LCD_RSTN_s1_address -> LT24_LCD_RSTN:address
	wire         mm_interconnect_0_lt24_lcd_rstn_s1_write;                     // mm_interconnect_0:LT24_LCD_RSTN_s1_write -> LT24_LCD_RSTN:write_n
	wire  [31:0] mm_interconnect_0_lt24_lcd_rstn_s1_writedata;                 // mm_interconnect_0:LT24_LCD_RSTN_s1_writedata -> LT24_LCD_RSTN:writedata
	wire         mm_interconnect_0_lt24_touch_penirq_n_s1_chipselect;          // mm_interconnect_0:LT24_TOUCH_PENIRQ_N_s1_chipselect -> LT24_TOUCH_PENIRQ_N:chipselect
	wire  [31:0] mm_interconnect_0_lt24_touch_penirq_n_s1_readdata;            // LT24_TOUCH_PENIRQ_N:readdata -> mm_interconnect_0:LT24_TOUCH_PENIRQ_N_s1_readdata
	wire   [1:0] mm_interconnect_0_lt24_touch_penirq_n_s1_address;             // mm_interconnect_0:LT24_TOUCH_PENIRQ_N_s1_address -> LT24_TOUCH_PENIRQ_N:address
	wire         mm_interconnect_0_lt24_touch_penirq_n_s1_write;               // mm_interconnect_0:LT24_TOUCH_PENIRQ_N_s1_write -> LT24_TOUCH_PENIRQ_N:write_n
	wire  [31:0] mm_interconnect_0_lt24_touch_penirq_n_s1_writedata;           // mm_interconnect_0:LT24_TOUCH_PENIRQ_N_s1_writedata -> LT24_TOUCH_PENIRQ_N:writedata
	wire  [31:0] mm_interconnect_0_lt24_touch_busy_s1_readdata;                // LT24_TOUCH_BUSY:readdata -> mm_interconnect_0:LT24_TOUCH_BUSY_s1_readdata
	wire   [1:0] mm_interconnect_0_lt24_touch_busy_s1_address;                 // mm_interconnect_0:LT24_TOUCH_BUSY_s1_address -> LT24_TOUCH_BUSY:address
	wire         mm_interconnect_0_pic_mem_s1_chipselect;                      // mm_interconnect_0:pic_mem_s1_chipselect -> pic_mem:chipselect
	wire  [15:0] mm_interconnect_0_pic_mem_s1_readdata;                        // pic_mem:readdata -> mm_interconnect_0:pic_mem_s1_readdata
	wire  [12:0] mm_interconnect_0_pic_mem_s1_address;                         // mm_interconnect_0:pic_mem_s1_address -> pic_mem:address
	wire   [1:0] mm_interconnect_0_pic_mem_s1_byteenable;                      // mm_interconnect_0:pic_mem_s1_byteenable -> pic_mem:byteenable
	wire         mm_interconnect_0_pic_mem_s1_write;                           // mm_interconnect_0:pic_mem_s1_write -> pic_mem:write
	wire  [15:0] mm_interconnect_0_pic_mem_s1_writedata;                       // mm_interconnect_0:pic_mem_s1_writedata -> pic_mem:writedata
	wire         mm_interconnect_0_pic_mem_s1_clken;                           // mm_interconnect_0:pic_mem_s1_clken -> pic_mem:clken
	wire         mm_interconnect_0_lt24_buffer_flag_s1_chipselect;             // mm_interconnect_0:LT24_buffer_flag_s1_chipselect -> LT24_buffer_flag:chipselect
	wire  [31:0] mm_interconnect_0_lt24_buffer_flag_s1_readdata;               // LT24_buffer_flag:readdata -> mm_interconnect_0:LT24_buffer_flag_s1_readdata
	wire   [1:0] mm_interconnect_0_lt24_buffer_flag_s1_address;                // mm_interconnect_0:LT24_buffer_flag_s1_address -> LT24_buffer_flag:address
	wire         mm_interconnect_0_lt24_buffer_flag_s1_write;                  // mm_interconnect_0:LT24_buffer_flag_s1_write -> LT24_buffer_flag:write_n
	wire  [31:0] mm_interconnect_0_lt24_buffer_flag_s1_writedata;              // mm_interconnect_0:LT24_buffer_flag_s1_writedata -> LT24_buffer_flag:writedata
	wire         mm_interconnect_0_background_mem_s1_chipselect;               // mm_interconnect_0:background_mem_s1_chipselect -> background_mem:chipselect
	wire  [15:0] mm_interconnect_0_background_mem_s1_readdata;                 // background_mem:readdata -> mm_interconnect_0:background_mem_s1_readdata
	wire  [12:0] mm_interconnect_0_background_mem_s1_address;                  // mm_interconnect_0:background_mem_s1_address -> background_mem:address
	wire   [1:0] mm_interconnect_0_background_mem_s1_byteenable;               // mm_interconnect_0:background_mem_s1_byteenable -> background_mem:byteenable
	wire         mm_interconnect_0_background_mem_s1_write;                    // mm_interconnect_0:background_mem_s1_write -> background_mem:write
	wire  [15:0] mm_interconnect_0_background_mem_s1_writedata;                // mm_interconnect_0:background_mem_s1_writedata -> background_mem:writedata
	wire         mm_interconnect_0_background_mem_s1_clken;                    // mm_interconnect_0:background_mem_s1_clken -> background_mem:clken
	wire  [31:0] mm_interconnect_0_gsensor_int_s1_readdata;                    // gsensor_int:readdata -> mm_interconnect_0:gsensor_int_s1_readdata
	wire   [1:0] mm_interconnect_0_gsensor_int_s1_address;                     // mm_interconnect_0:gsensor_int_s1_address -> gsensor_int:address
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;                // mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;                  // sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                   // mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                     // mm_interconnect_0:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;                 // mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_0_sdram_controler_s1_chipselect;              // mm_interconnect_0:SDRAM_Controler_s1_chipselect -> SDRAM_Controler:az_cs
	wire  [15:0] mm_interconnect_0_sdram_controler_s1_readdata;                // SDRAM_Controler:za_data -> mm_interconnect_0:SDRAM_Controler_s1_readdata
	wire         mm_interconnect_0_sdram_controler_s1_waitrequest;             // SDRAM_Controler:za_waitrequest -> mm_interconnect_0:SDRAM_Controler_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_controler_s1_address;                 // mm_interconnect_0:SDRAM_Controler_s1_address -> SDRAM_Controler:az_addr
	wire         mm_interconnect_0_sdram_controler_s1_read;                    // mm_interconnect_0:SDRAM_Controler_s1_read -> SDRAM_Controler:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_controler_s1_byteenable;              // mm_interconnect_0:SDRAM_Controler_s1_byteenable -> SDRAM_Controler:az_be_n
	wire         mm_interconnect_0_sdram_controler_s1_readdatavalid;           // SDRAM_Controler:za_valid -> mm_interconnect_0:SDRAM_Controler_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controler_s1_write;                   // mm_interconnect_0:SDRAM_Controler_s1_write -> SDRAM_Controler:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_controler_s1_writedata;               // mm_interconnect_0:SDRAM_Controler_s1_writedata -> SDRAM_Controler:az_data
	wire         mm_interconnect_0_timer_timestamp_s1_chipselect;              // mm_interconnect_0:timer_timestamp_s1_chipselect -> timer_timestamp:chipselect
	wire  [15:0] mm_interconnect_0_timer_timestamp_s1_readdata;                // timer_timestamp:readdata -> mm_interconnect_0:timer_timestamp_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_timestamp_s1_address;                 // mm_interconnect_0:timer_timestamp_s1_address -> timer_timestamp:address
	wire         mm_interconnect_0_timer_timestamp_s1_write;                   // mm_interconnect_0:timer_timestamp_s1_write -> timer_timestamp:write_n
	wire  [15:0] mm_interconnect_0_timer_timestamp_s1_writedata;               // mm_interconnect_0:timer_timestamp_s1_writedata -> timer_timestamp:writedata
	wire         mm_interconnect_0_gsensor_spi_slave_chipselect;               // mm_interconnect_0:gsensor_spi_slave_chipselect -> gsensor_spi:s_chipselect
	wire   [7:0] mm_interconnect_0_gsensor_spi_slave_readdata;                 // gsensor_spi:s_readdata -> mm_interconnect_0:gsensor_spi_slave_readdata
	wire   [3:0] mm_interconnect_0_gsensor_spi_slave_address;                  // mm_interconnect_0:gsensor_spi_slave_address -> gsensor_spi:s_address
	wire         mm_interconnect_0_gsensor_spi_slave_read;                     // mm_interconnect_0:gsensor_spi_slave_read -> gsensor_spi:s_read
	wire         mm_interconnect_0_gsensor_spi_slave_write;                    // mm_interconnect_0:gsensor_spi_slave_write -> gsensor_spi:s_write
	wire   [7:0] mm_interconnect_0_gsensor_spi_slave_writedata;                // mm_interconnect_0:gsensor_spi_slave_writedata -> gsensor_spi:s_writedata
	wire         mm_interconnect_0_lt24_touch_spi_spi_control_port_chipselect; // mm_interconnect_0:LT24_TOUCH_SPI_spi_control_port_chipselect -> LT24_TOUCH_SPI:spi_select
	wire  [15:0] mm_interconnect_0_lt24_touch_spi_spi_control_port_readdata;   // LT24_TOUCH_SPI:data_to_cpu -> mm_interconnect_0:LT24_TOUCH_SPI_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_lt24_touch_spi_spi_control_port_address;    // mm_interconnect_0:LT24_TOUCH_SPI_spi_control_port_address -> LT24_TOUCH_SPI:mem_addr
	wire         mm_interconnect_0_lt24_touch_spi_spi_control_port_read;       // mm_interconnect_0:LT24_TOUCH_SPI_spi_control_port_read -> LT24_TOUCH_SPI:read_n
	wire         mm_interconnect_0_lt24_touch_spi_spi_control_port_write;      // mm_interconnect_0:LT24_TOUCH_SPI_spi_control_port_write -> LT24_TOUCH_SPI:write_n
	wire  [15:0] mm_interconnect_0_lt24_touch_spi_spi_control_port_writedata;  // mm_interconnect_0:LT24_TOUCH_SPI_spi_control_port_writedata -> LT24_TOUCH_SPI:data_from_cpu
	wire         irq_mapper_receiver2_irq;                                     // JTAG_UART:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver4_irq;                                     // LT24_TOUCH_SPI:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                     // LT24_TOUCH_PENIRQ_N:irq -> irq_mapper:receiver5_irq
	wire  [31:0] cpu_d_irq_irq;                                                // irq_mapper:sender_irq -> CPU:d_irq
	wire         irq_mapper_receiver0_irq;                                     // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                // cycloneSPI:ins_irq0_irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                     // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                            // LT24_interface_irq_0:ins_irq0_irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver3_irq;                                     // irq_synchronizer_002:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                            // TIMER:irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver6_irq;                                     // irq_synchronizer_003:sender_irq -> irq_mapper:receiver6_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                            // sys_clk_timer:irq -> irq_synchronizer_003:receiver_irq
	wire         irq_mapper_receiver7_irq;                                     // irq_synchronizer_004:sender_irq -> irq_mapper:receiver7_irq
	wire   [0:0] irq_synchronizer_004_receiver_irq;                            // timer_timestamp:irq -> irq_synchronizer_004:receiver_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [ALT_PLL:reset, background_mem:reset, background_mem:reset2, mm_interconnect_0:ALT_PLL_inclk_interface_reset_reset_bridge_in_reset_reset, pic_mem:reset, pic_mem:reset2]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [background_mem:reset_req, background_mem:reset_req2, pic_mem:reset_req, pic_mem:reset_req2, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                            // CPU:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [CPU:reset_n, JTAG_UART:rst_n, LT24_CTRL:reset_n, LT24_LCD_RSTN:reset_n, LT24_TOUCH_BUSY:reset_n, LT24_TOUCH_PENIRQ_N:reset_n, LT24_TOUCH_SPI:reset_n, SDRAM_Controler:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, mm_interconnect_0:CPU_reset_n_reset_bridge_in_reset_reset, rst_translator_001:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                       // rst_controller_001:reset_req -> [CPU:reset_req, rst_translator_001:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                           // rst_controller_002:reset_out -> [KEY:reset_n, LED_CTRL:RST, TIMER:reset_n, irq_synchronizer_002:receiver_reset, mm_interconnect_0:LED_CTRL_reset_sink_reset_bridge_in_reset_reset]
	wire         rst_controller_003_reset_out_reset;                           // rst_controller_003:reset_out -> [LT24_buffer_flag:reset_n, LT24_interface_irq_0:reset_reset, gsensor_int:reset_n, gsensor_spi:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, mm_interconnect_0:LT24_interface_irq_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:cycloneSPI_reset_sink_reset_bridge_in_reset_reset, sys_clk_timer:reset_n, timer_timestamp:reset_n]

	DE0_LT24_SOPC_ALT_PLL alt_pll (
		.clk       (clk_clk),                                       //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                // inclk_interface_reset.reset
		.read      (mm_interconnect_0_alt_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_alt_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_alt_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_alt_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_alt_pll_pll_slave_writedata), //                      .writedata
		.c0        (alt_pll_c0_clk),                                //                    c0.clk
		.c1        (alt_pll_c1_clk),                                //                    c1.clk
		.c2        (alt_pll_c2_clk),                                //                    c2.clk
		.c3        (alt_pll_c3_clk),                                //                    c3.clk
		.c4        (),                                              //                    c4.clk
		.areset    (alt_pll_areset_conduit_export),                 //        areset_conduit.export
		.locked    (alt_pll_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (alt_pll_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	DE0_LT24_SOPC_CPU cpu (
		.clk                                   (alt_pll_c0_clk),                                      //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	DE0_LT24_SOPC_JTAG_UART jtag_uart (
		.clk            (alt_pll_c0_clk),                                            //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	DE0_LT24_SOPC_KEY key (
		.clk      (alt_pll_c2_clk),                      //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_key_s1_address),    //                  s1.address
		.readdata (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port  (from_key_export)                      // external_connection.export
	);

	LED_Controller led_ctrl (
		.CLK   (alt_pll_c2_clk),                                      //          clock.clk
		.WRITE (mm_interconnect_0_led_ctrl_avalon_slave_0_write),     // avalon_slave_0.write
		.READ  (mm_interconnect_0_led_ctrl_avalon_slave_0_read),      //               .read
		.ADDR  (mm_interconnect_0_led_ctrl_avalon_slave_0_address),   //               .address
		.WDATA (mm_interconnect_0_led_ctrl_avalon_slave_0_writedata), //               .writedata
		.RDATA (mm_interconnect_0_led_ctrl_avalon_slave_0_readdata),  //               .readdata
		.RST   (rst_controller_002_reset_out_reset),                  //     reset_sink.reset
		.LED   (to_led_export)                                        //    conduit_end.export
	);

	LT24_Controller lt24_ctrl (
		.clk            (alt_pll_c0_clk),                                         //          clock.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                    //          reset.reset_n
		.s_chipselect_n (~mm_interconnect_0_lt24_ctrl_avalon_slave_0_chipselect), // avalon_slave_0.chipselect_n
		.s_write_n      (~mm_interconnect_0_lt24_ctrl_avalon_slave_0_write),      //               .write_n
		.s_writedata    (mm_interconnect_0_lt24_ctrl_avalon_slave_0_writedata),   //               .writedata
		.s_address      (mm_interconnect_0_lt24_ctrl_avalon_slave_0_address),     //               .address
		.lt24_cs        (lt24_conduit_cs),                                        //    conduit_end.export
		.lt24_rs        (lt24_conduit_rs),                                        //               .export
		.lt24_rd        (lt24_conduit_rd),                                        //               .export
		.lt24_wr        (lt24_conduit_wr),                                        //               .export
		.lt24_data      (lt24_conduit_data)                                       //               .export
	);

	DE0_LT24_SOPC_LT24_LCD_RSTN lt24_lcd_rstn (
		.clk        (alt_pll_c0_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_lt24_lcd_rstn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lt24_lcd_rstn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lt24_lcd_rstn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lt24_lcd_rstn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lt24_lcd_rstn_s1_readdata),   //                    .readdata
		.out_port   (lt24_lcd_rstn_export)                           // external_connection.export
	);

	DE0_LT24_SOPC_LT24_TOUCH_BUSY lt24_touch_busy (
		.clk      (alt_pll_c0_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_lt24_touch_busy_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_lt24_touch_busy_s1_readdata), //                    .readdata
		.in_port  (lt24_touch_busy_export)                         // external_connection.export
	);

	DE0_LT24_SOPC_LT24_TOUCH_PENIRQ_N lt24_touch_penirq_n (
		.clk        (alt_pll_c0_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_lt24_touch_penirq_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lt24_touch_penirq_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lt24_touch_penirq_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lt24_touch_penirq_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lt24_touch_penirq_n_s1_readdata),   //                    .readdata
		.in_port    (lt24_touch_penirq_n_export),                          // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                             //                 irq.irq
	);

	DE0_LT24_SOPC_LT24_TOUCH_SPI lt24_touch_spi (
		.clk           (alt_pll_c0_clk),                                               //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                          //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_lt24_touch_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_lt24_touch_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_lt24_touch_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_lt24_touch_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_lt24_touch_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_lt24_touch_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver4_irq),                                     //              irq.irq
		.MISO          (lt24_touch_spi_MISO),                                          //         external.export
		.MOSI          (lt24_touch_spi_MOSI),                                          //                 .export
		.SCLK          (lt24_touch_spi_SCLK),                                          //                 .export
		.SS_n          (lt24_touch_spi_SS_n)                                           //                 .export
	);

	DE0_LT24_SOPC_LT24_LCD_RSTN lt24_buffer_flag (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_lt24_buffer_flag_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lt24_buffer_flag_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lt24_buffer_flag_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lt24_buffer_flag_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lt24_buffer_flag_s1_readdata),   //                    .readdata
		.out_port   (lt24_buffer_flag_external_connection_export)       // external_connection.export
	);

	LT24_interface_irq lt24_interface_irq_0 (
		.avs_s0_address     (mm_interconnect_0_lt24_interface_irq_0_avs_s0_address),     //      avs_s0.address
		.avs_s0_read        (mm_interconnect_0_lt24_interface_irq_0_avs_s0_read),        //            .read
		.avs_s0_readdata    (mm_interconnect_0_lt24_interface_irq_0_avs_s0_readdata),    //            .readdata
		.avs_s0_write       (mm_interconnect_0_lt24_interface_irq_0_avs_s0_write),       //            .write
		.avs_s0_writedata   (mm_interconnect_0_lt24_interface_irq_0_avs_s0_writedata),   //            .writedata
		.avs_s0_waitrequest (mm_interconnect_0_lt24_interface_irq_0_avs_s0_waitrequest), //            .waitrequest
		.clock_clk          (clk_clk),                                                   //       clock.clk
		.reset_reset        (rst_controller_003_reset_out_reset),                        //       reset.reset
		.ins_irq0_irq       (irq_synchronizer_001_receiver_irq),                         //    ins_irq0.irq
		.finish_flag        (lt24_conduit_0_finish_flag),                                // conduit_end.finish_flag
		.counter            (lt24_conduit_0_counter),                                    //            .counter
		.pattern            (lt24_conduit_0_pattern),                                    //            .pattern
		.vx                 (lt24_conduit_0_vx),                                         //            .vx
		.vy                 (lt24_conduit_0_vy),                                         //            .vy
		.lt24_coin_x0       (lt24_conduit_0_lt24_coin_x0),                               //            .lt24_coin_x0
		.lt24_coin_y0       (lt24_conduit_0_lt42_coin_y0),                               //            .lt42_coin_y0
		.lt24_coin_x        (lt24_conduit_0_lt24_coinx),                                 //            .lt24_coinx
		.lt24_coin_y        (lt24_conduit_0_lt24_coin_y),                                //            .lt24_coin_y
		.lt24_coin_vx0      (lt24_conduit_0_lt24_coin_vx0),                              //            .lt24_coin_vx0
		.lt24_coin_vy0      (lt24_conduit_0_lt24_coin_vy0)                               //            .lt24_coin_vy0
	);

	DE0_LT24_SOPC_SDRAM_Controler sdram_controler (
		.clk            (alt_pll_c0_clk),                                     //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controler_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controler_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controler_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controler_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controler_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controler_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controler_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controler_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controler_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controler_wire_addr),                          //  wire.export
		.zs_ba          (sdram_controler_wire_ba),                            //      .export
		.zs_cas_n       (sdram_controler_wire_cas_n),                         //      .export
		.zs_cke         (sdram_controler_wire_cke),                           //      .export
		.zs_cs_n        (sdram_controler_wire_cs_n),                          //      .export
		.zs_dq          (sdram_controler_wire_dq),                            //      .export
		.zs_dqm         (sdram_controler_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_controler_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_controler_wire_we_n)                           //      .export
	);

	DE0_LT24_SOPC_TIMER timer (
		.clk        (alt_pll_c2_clk),                        //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_002_receiver_irq)      //   irq.irq
	);

	DE0_LT24_SOPC_background_mem background_mem (
		.clk         (clk_clk),                                        //   clk1.clk
		.address     (mm_interconnect_0_background_mem_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_background_mem_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_background_mem_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_background_mem_s1_write),      //       .write
		.readdata    (mm_interconnect_0_background_mem_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_background_mem_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_background_mem_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),             //       .reset_req
		.address2    (background_mem_s2_address),                      //     s2.address
		.chipselect2 (background_mem_s2_chipselect),                   //       .chipselect
		.clken2      (background_mem_s2_clken),                        //       .clken
		.write2      (background_mem_s2_write),                        //       .write
		.readdata2   (background_mem_s2_readdata),                     //       .readdata
		.writedata2  (background_mem_s2_writedata),                    //       .writedata
		.byteenable2 (background_mem_s2_byteenable),                   //       .byteenable
		.clk2        (clk_clk),                                        //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                 // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req)              //       .reset_req
	);

	MyCycloneSPI cyclonespi (
		.clk                (clk_clk),                                         //    clock_sink.clk
		.reset              (~reset_reset_n),                                  //    reset_sink.reset
		.SPI_clk            (cyclonespi_spi_interface_SPI_clk),                // SPI_interface.SPI_clk
		.SPI_CS             (cyclonespi_spi_interface_SPI_CS),                 //              .SPI_CS
		.SPI_SDI            (cyclonespi_spi_interface_SPI_SDI),                //              .SPI_SDI
		.SPI_SDO            (cyclonespi_spi_interface_SPI_SDO),                //              .SPI_SDO
		.data_out           (cyclonespi_spi_interface_data_out),               //              .data_out
		.data_out_enable    (cyclonespi_spi_interface_data_out_enable),        //              .data_out_enable
		.Config             (cyclonespi_spi_interface_config),                 //              .config
		.spi_irq            (cyclonespi_spi_interface_spi_irq),                //              .spi_irq
		.avs_s0_address     (mm_interconnect_0_cyclonespi_avs_s0_address),     //        avs_s0.address
		.avs_s0_read        (mm_interconnect_0_cyclonespi_avs_s0_read),        //              .read
		.avs_s0_readdata    (mm_interconnect_0_cyclonespi_avs_s0_readdata),    //              .readdata
		.avs_s0_write       (mm_interconnect_0_cyclonespi_avs_s0_write),       //              .write
		.avs_s0_writedata   (mm_interconnect_0_cyclonespi_avs_s0_writedata),   //              .writedata
		.avs_s0_waitrequest (mm_interconnect_0_cyclonespi_avs_s0_waitrequest), //              .waitrequest
		.ins_irq0_irq       (irq_synchronizer_receiver_irq)                    //      ins_irq0.irq
	);

	DE0_LT24_SOPC_LT24_TOUCH_BUSY gsensor_int (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_gsensor_int_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_gsensor_int_s1_readdata), //                    .readdata
		.in_port  (gsensor_int_external_connection_export)     // external_connection.export
	);

	TERASIC_SPI_3WIRE gsensor_spi (
		.clk          (clk_clk),                                        //       clock_reset.clk
		.reset_n      (~rst_controller_003_reset_out_reset),            // clock_reset_reset.reset_n
		.s_chipselect (mm_interconnect_0_gsensor_spi_slave_chipselect), //             slave.chipselect
		.s_address    (mm_interconnect_0_gsensor_spi_slave_address),    //                  .address
		.s_write      (mm_interconnect_0_gsensor_spi_slave_write),      //                  .write
		.s_writedata  (mm_interconnect_0_gsensor_spi_slave_writedata),  //                  .writedata
		.s_read       (mm_interconnect_0_gsensor_spi_slave_read),       //                  .read
		.s_readdata   (mm_interconnect_0_gsensor_spi_slave_readdata),   //                  .readdata
		.SPI_SDIO     (gsensor_spi_conduit_end_SDIO),                   //       conduit_end.export
		.SPI_SCLK     (gsensor_spi_conduit_end_SCLK),                   //                  .export
		.SPI_CS_n     (gsensor_spi_conduit_end_CS_n)                    //                  .export
	);

	DE0_LT24_SOPC_pic_mem pic_mem (
		.clk         (clk_clk),                                 //   clk1.clk
		.address     (mm_interconnect_0_pic_mem_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_pic_mem_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_pic_mem_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_pic_mem_s1_write),      //       .write
		.readdata    (mm_interconnect_0_pic_mem_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_pic_mem_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_pic_mem_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),      //       .reset_req
		.address2    (pic_mem_s2_address),                      //     s2.address
		.chipselect2 (pic_mem_s2_chipselect),                   //       .chipselect
		.clken2      (pic_mem_s2_clken),                        //       .clken
		.write2      (pic_mem_s2_write),                        //       .write
		.readdata2   (pic_mem_s2_readdata),                     //       .readdata
		.writedata2  (pic_mem_s2_writedata),                    //       .writedata
		.byteenable2 (pic_mem_s2_byteenable),                   //       .byteenable
		.clk2        (clk_clk),                                 //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),          // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req)       //       .reset_req
	);

	DE0_LT24_SOPC_sys_clk_timer sys_clk_timer (
		.clk        (clk_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_003_receiver_irq)              //   irq.irq
	);

	DE0_LT24_SOPC_sys_clk_timer timer_timestamp (
		.clk        (clk_clk),                                         //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),             // reset.reset_n
		.address    (mm_interconnect_0_timer_timestamp_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_timestamp_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_timestamp_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_timestamp_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_timestamp_s1_write),     //      .write_n
		.irq        (irq_synchronizer_004_receiver_irq)                //   irq.irq
	);

	DE0_LT24_SOPC_mm_interconnect_0 mm_interconnect_0 (
		.ALT_PLL_c0_clk                                            (alt_pll_c0_clk),                                               //                                          ALT_PLL_c0.clk
		.ALT_PLL_c2_clk                                            (alt_pll_c2_clk),                                               //                                          ALT_PLL_c2.clk
		.CLK_50_clk_clk                                            (clk_clk),                                                      //                                          CLK_50_clk.clk
		.ALT_PLL_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // ALT_PLL_inclk_interface_reset_reset_bridge_in_reset.reset
		.CPU_reset_n_reset_bridge_in_reset_reset                   (rst_controller_001_reset_out_reset),                           //                   CPU_reset_n_reset_bridge_in_reset.reset
		.cycloneSPI_reset_sink_reset_bridge_in_reset_reset         (rst_controller_003_reset_out_reset),                           //         cycloneSPI_reset_sink_reset_bridge_in_reset.reset
		.LED_CTRL_reset_sink_reset_bridge_in_reset_reset           (rst_controller_002_reset_out_reset),                           //           LED_CTRL_reset_sink_reset_bridge_in_reset.reset
		.LT24_interface_irq_0_reset_reset_bridge_in_reset_reset    (rst_controller_003_reset_out_reset),                           //    LT24_interface_irq_0_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address                                   (cpu_data_master_address),                                      //                                     CPU_data_master.address
		.CPU_data_master_waitrequest                               (cpu_data_master_waitrequest),                                  //                                                    .waitrequest
		.CPU_data_master_byteenable                                (cpu_data_master_byteenable),                                   //                                                    .byteenable
		.CPU_data_master_read                                      (cpu_data_master_read),                                         //                                                    .read
		.CPU_data_master_readdata                                  (cpu_data_master_readdata),                                     //                                                    .readdata
		.CPU_data_master_readdatavalid                             (cpu_data_master_readdatavalid),                                //                                                    .readdatavalid
		.CPU_data_master_write                                     (cpu_data_master_write),                                        //                                                    .write
		.CPU_data_master_writedata                                 (cpu_data_master_writedata),                                    //                                                    .writedata
		.CPU_data_master_debugaccess                               (cpu_data_master_debugaccess),                                  //                                                    .debugaccess
		.CPU_instruction_master_address                            (cpu_instruction_master_address),                               //                              CPU_instruction_master.address
		.CPU_instruction_master_waitrequest                        (cpu_instruction_master_waitrequest),                           //                                                    .waitrequest
		.CPU_instruction_master_read                               (cpu_instruction_master_read),                                  //                                                    .read
		.CPU_instruction_master_readdata                           (cpu_instruction_master_readdata),                              //                                                    .readdata
		.CPU_instruction_master_readdatavalid                      (cpu_instruction_master_readdatavalid),                         //                                                    .readdatavalid
		.ALT_PLL_pll_slave_address                                 (mm_interconnect_0_alt_pll_pll_slave_address),                  //                                   ALT_PLL_pll_slave.address
		.ALT_PLL_pll_slave_write                                   (mm_interconnect_0_alt_pll_pll_slave_write),                    //                                                    .write
		.ALT_PLL_pll_slave_read                                    (mm_interconnect_0_alt_pll_pll_slave_read),                     //                                                    .read
		.ALT_PLL_pll_slave_readdata                                (mm_interconnect_0_alt_pll_pll_slave_readdata),                 //                                                    .readdata
		.ALT_PLL_pll_slave_writedata                               (mm_interconnect_0_alt_pll_pll_slave_writedata),                //                                                    .writedata
		.background_mem_s1_address                                 (mm_interconnect_0_background_mem_s1_address),                  //                                   background_mem_s1.address
		.background_mem_s1_write                                   (mm_interconnect_0_background_mem_s1_write),                    //                                                    .write
		.background_mem_s1_readdata                                (mm_interconnect_0_background_mem_s1_readdata),                 //                                                    .readdata
		.background_mem_s1_writedata                               (mm_interconnect_0_background_mem_s1_writedata),                //                                                    .writedata
		.background_mem_s1_byteenable                              (mm_interconnect_0_background_mem_s1_byteenable),               //                                                    .byteenable
		.background_mem_s1_chipselect                              (mm_interconnect_0_background_mem_s1_chipselect),               //                                                    .chipselect
		.background_mem_s1_clken                                   (mm_interconnect_0_background_mem_s1_clken),                    //                                                    .clken
		.CPU_jtag_debug_module_address                             (mm_interconnect_0_cpu_jtag_debug_module_address),              //                               CPU_jtag_debug_module.address
		.CPU_jtag_debug_module_write                               (mm_interconnect_0_cpu_jtag_debug_module_write),                //                                                    .write
		.CPU_jtag_debug_module_read                                (mm_interconnect_0_cpu_jtag_debug_module_read),                 //                                                    .read
		.CPU_jtag_debug_module_readdata                            (mm_interconnect_0_cpu_jtag_debug_module_readdata),             //                                                    .readdata
		.CPU_jtag_debug_module_writedata                           (mm_interconnect_0_cpu_jtag_debug_module_writedata),            //                                                    .writedata
		.CPU_jtag_debug_module_byteenable                          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),           //                                                    .byteenable
		.CPU_jtag_debug_module_waitrequest                         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),          //                                                    .waitrequest
		.CPU_jtag_debug_module_debugaccess                         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),          //                                                    .debugaccess
		.cycloneSPI_avs_s0_address                                 (mm_interconnect_0_cyclonespi_avs_s0_address),                  //                                   cycloneSPI_avs_s0.address
		.cycloneSPI_avs_s0_write                                   (mm_interconnect_0_cyclonespi_avs_s0_write),                    //                                                    .write
		.cycloneSPI_avs_s0_read                                    (mm_interconnect_0_cyclonespi_avs_s0_read),                     //                                                    .read
		.cycloneSPI_avs_s0_readdata                                (mm_interconnect_0_cyclonespi_avs_s0_readdata),                 //                                                    .readdata
		.cycloneSPI_avs_s0_writedata                               (mm_interconnect_0_cyclonespi_avs_s0_writedata),                //                                                    .writedata
		.cycloneSPI_avs_s0_waitrequest                             (mm_interconnect_0_cyclonespi_avs_s0_waitrequest),              //                                                    .waitrequest
		.gsensor_int_s1_address                                    (mm_interconnect_0_gsensor_int_s1_address),                     //                                      gsensor_int_s1.address
		.gsensor_int_s1_readdata                                   (mm_interconnect_0_gsensor_int_s1_readdata),                    //                                                    .readdata
		.gsensor_spi_slave_address                                 (mm_interconnect_0_gsensor_spi_slave_address),                  //                                   gsensor_spi_slave.address
		.gsensor_spi_slave_write                                   (mm_interconnect_0_gsensor_spi_slave_write),                    //                                                    .write
		.gsensor_spi_slave_read                                    (mm_interconnect_0_gsensor_spi_slave_read),                     //                                                    .read
		.gsensor_spi_slave_readdata                                (mm_interconnect_0_gsensor_spi_slave_readdata),                 //                                                    .readdata
		.gsensor_spi_slave_writedata                               (mm_interconnect_0_gsensor_spi_slave_writedata),                //                                                    .writedata
		.gsensor_spi_slave_chipselect                              (mm_interconnect_0_gsensor_spi_slave_chipselect),               //                                                    .chipselect
		.JTAG_UART_avalon_jtag_slave_address                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),        //                         JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),          //                                                    .write
		.JTAG_UART_avalon_jtag_slave_read                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),           //                                                    .read
		.JTAG_UART_avalon_jtag_slave_readdata                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),       //                                                    .readdata
		.JTAG_UART_avalon_jtag_slave_writedata                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),      //                                                    .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),    //                                                    .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),     //                                                    .chipselect
		.KEY_s1_address                                            (mm_interconnect_0_key_s1_address),                             //                                              KEY_s1.address
		.KEY_s1_readdata                                           (mm_interconnect_0_key_s1_readdata),                            //                                                    .readdata
		.LED_CTRL_avalon_slave_0_address                           (mm_interconnect_0_led_ctrl_avalon_slave_0_address),            //                             LED_CTRL_avalon_slave_0.address
		.LED_CTRL_avalon_slave_0_write                             (mm_interconnect_0_led_ctrl_avalon_slave_0_write),              //                                                    .write
		.LED_CTRL_avalon_slave_0_read                              (mm_interconnect_0_led_ctrl_avalon_slave_0_read),               //                                                    .read
		.LED_CTRL_avalon_slave_0_readdata                          (mm_interconnect_0_led_ctrl_avalon_slave_0_readdata),           //                                                    .readdata
		.LED_CTRL_avalon_slave_0_writedata                         (mm_interconnect_0_led_ctrl_avalon_slave_0_writedata),          //                                                    .writedata
		.LT24_buffer_flag_s1_address                               (mm_interconnect_0_lt24_buffer_flag_s1_address),                //                                 LT24_buffer_flag_s1.address
		.LT24_buffer_flag_s1_write                                 (mm_interconnect_0_lt24_buffer_flag_s1_write),                  //                                                    .write
		.LT24_buffer_flag_s1_readdata                              (mm_interconnect_0_lt24_buffer_flag_s1_readdata),               //                                                    .readdata
		.LT24_buffer_flag_s1_writedata                             (mm_interconnect_0_lt24_buffer_flag_s1_writedata),              //                                                    .writedata
		.LT24_buffer_flag_s1_chipselect                            (mm_interconnect_0_lt24_buffer_flag_s1_chipselect),             //                                                    .chipselect
		.LT24_CTRL_avalon_slave_0_address                          (mm_interconnect_0_lt24_ctrl_avalon_slave_0_address),           //                            LT24_CTRL_avalon_slave_0.address
		.LT24_CTRL_avalon_slave_0_write                            (mm_interconnect_0_lt24_ctrl_avalon_slave_0_write),             //                                                    .write
		.LT24_CTRL_avalon_slave_0_writedata                        (mm_interconnect_0_lt24_ctrl_avalon_slave_0_writedata),         //                                                    .writedata
		.LT24_CTRL_avalon_slave_0_chipselect                       (mm_interconnect_0_lt24_ctrl_avalon_slave_0_chipselect),        //                                                    .chipselect
		.LT24_interface_irq_0_avs_s0_address                       (mm_interconnect_0_lt24_interface_irq_0_avs_s0_address),        //                         LT24_interface_irq_0_avs_s0.address
		.LT24_interface_irq_0_avs_s0_write                         (mm_interconnect_0_lt24_interface_irq_0_avs_s0_write),          //                                                    .write
		.LT24_interface_irq_0_avs_s0_read                          (mm_interconnect_0_lt24_interface_irq_0_avs_s0_read),           //                                                    .read
		.LT24_interface_irq_0_avs_s0_readdata                      (mm_interconnect_0_lt24_interface_irq_0_avs_s0_readdata),       //                                                    .readdata
		.LT24_interface_irq_0_avs_s0_writedata                     (mm_interconnect_0_lt24_interface_irq_0_avs_s0_writedata),      //                                                    .writedata
		.LT24_interface_irq_0_avs_s0_waitrequest                   (mm_interconnect_0_lt24_interface_irq_0_avs_s0_waitrequest),    //                                                    .waitrequest
		.LT24_LCD_RSTN_s1_address                                  (mm_interconnect_0_lt24_lcd_rstn_s1_address),                   //                                    LT24_LCD_RSTN_s1.address
		.LT24_LCD_RSTN_s1_write                                    (mm_interconnect_0_lt24_lcd_rstn_s1_write),                     //                                                    .write
		.LT24_LCD_RSTN_s1_readdata                                 (mm_interconnect_0_lt24_lcd_rstn_s1_readdata),                  //                                                    .readdata
		.LT24_LCD_RSTN_s1_writedata                                (mm_interconnect_0_lt24_lcd_rstn_s1_writedata),                 //                                                    .writedata
		.LT24_LCD_RSTN_s1_chipselect                               (mm_interconnect_0_lt24_lcd_rstn_s1_chipselect),                //                                                    .chipselect
		.LT24_TOUCH_BUSY_s1_address                                (mm_interconnect_0_lt24_touch_busy_s1_address),                 //                                  LT24_TOUCH_BUSY_s1.address
		.LT24_TOUCH_BUSY_s1_readdata                               (mm_interconnect_0_lt24_touch_busy_s1_readdata),                //                                                    .readdata
		.LT24_TOUCH_PENIRQ_N_s1_address                            (mm_interconnect_0_lt24_touch_penirq_n_s1_address),             //                              LT24_TOUCH_PENIRQ_N_s1.address
		.LT24_TOUCH_PENIRQ_N_s1_write                              (mm_interconnect_0_lt24_touch_penirq_n_s1_write),               //                                                    .write
		.LT24_TOUCH_PENIRQ_N_s1_readdata                           (mm_interconnect_0_lt24_touch_penirq_n_s1_readdata),            //                                                    .readdata
		.LT24_TOUCH_PENIRQ_N_s1_writedata                          (mm_interconnect_0_lt24_touch_penirq_n_s1_writedata),           //                                                    .writedata
		.LT24_TOUCH_PENIRQ_N_s1_chipselect                         (mm_interconnect_0_lt24_touch_penirq_n_s1_chipselect),          //                                                    .chipselect
		.LT24_TOUCH_SPI_spi_control_port_address                   (mm_interconnect_0_lt24_touch_spi_spi_control_port_address),    //                     LT24_TOUCH_SPI_spi_control_port.address
		.LT24_TOUCH_SPI_spi_control_port_write                     (mm_interconnect_0_lt24_touch_spi_spi_control_port_write),      //                                                    .write
		.LT24_TOUCH_SPI_spi_control_port_read                      (mm_interconnect_0_lt24_touch_spi_spi_control_port_read),       //                                                    .read
		.LT24_TOUCH_SPI_spi_control_port_readdata                  (mm_interconnect_0_lt24_touch_spi_spi_control_port_readdata),   //                                                    .readdata
		.LT24_TOUCH_SPI_spi_control_port_writedata                 (mm_interconnect_0_lt24_touch_spi_spi_control_port_writedata),  //                                                    .writedata
		.LT24_TOUCH_SPI_spi_control_port_chipselect                (mm_interconnect_0_lt24_touch_spi_spi_control_port_chipselect), //                                                    .chipselect
		.pic_mem_s1_address                                        (mm_interconnect_0_pic_mem_s1_address),                         //                                          pic_mem_s1.address
		.pic_mem_s1_write                                          (mm_interconnect_0_pic_mem_s1_write),                           //                                                    .write
		.pic_mem_s1_readdata                                       (mm_interconnect_0_pic_mem_s1_readdata),                        //                                                    .readdata
		.pic_mem_s1_writedata                                      (mm_interconnect_0_pic_mem_s1_writedata),                       //                                                    .writedata
		.pic_mem_s1_byteenable                                     (mm_interconnect_0_pic_mem_s1_byteenable),                      //                                                    .byteenable
		.pic_mem_s1_chipselect                                     (mm_interconnect_0_pic_mem_s1_chipselect),                      //                                                    .chipselect
		.pic_mem_s1_clken                                          (mm_interconnect_0_pic_mem_s1_clken),                           //                                                    .clken
		.SDRAM_Controler_s1_address                                (mm_interconnect_0_sdram_controler_s1_address),                 //                                  SDRAM_Controler_s1.address
		.SDRAM_Controler_s1_write                                  (mm_interconnect_0_sdram_controler_s1_write),                   //                                                    .write
		.SDRAM_Controler_s1_read                                   (mm_interconnect_0_sdram_controler_s1_read),                    //                                                    .read
		.SDRAM_Controler_s1_readdata                               (mm_interconnect_0_sdram_controler_s1_readdata),                //                                                    .readdata
		.SDRAM_Controler_s1_writedata                              (mm_interconnect_0_sdram_controler_s1_writedata),               //                                                    .writedata
		.SDRAM_Controler_s1_byteenable                             (mm_interconnect_0_sdram_controler_s1_byteenable),              //                                                    .byteenable
		.SDRAM_Controler_s1_readdatavalid                          (mm_interconnect_0_sdram_controler_s1_readdatavalid),           //                                                    .readdatavalid
		.SDRAM_Controler_s1_waitrequest                            (mm_interconnect_0_sdram_controler_s1_waitrequest),             //                                                    .waitrequest
		.SDRAM_Controler_s1_chipselect                             (mm_interconnect_0_sdram_controler_s1_chipselect),              //                                                    .chipselect
		.sys_clk_timer_s1_address                                  (mm_interconnect_0_sys_clk_timer_s1_address),                   //                                    sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                                    (mm_interconnect_0_sys_clk_timer_s1_write),                     //                                                    .write
		.sys_clk_timer_s1_readdata                                 (mm_interconnect_0_sys_clk_timer_s1_readdata),                  //                                                    .readdata
		.sys_clk_timer_s1_writedata                                (mm_interconnect_0_sys_clk_timer_s1_writedata),                 //                                                    .writedata
		.sys_clk_timer_s1_chipselect                               (mm_interconnect_0_sys_clk_timer_s1_chipselect),                //                                                    .chipselect
		.TIMER_s1_address                                          (mm_interconnect_0_timer_s1_address),                           //                                            TIMER_s1.address
		.TIMER_s1_write                                            (mm_interconnect_0_timer_s1_write),                             //                                                    .write
		.TIMER_s1_readdata                                         (mm_interconnect_0_timer_s1_readdata),                          //                                                    .readdata
		.TIMER_s1_writedata                                        (mm_interconnect_0_timer_s1_writedata),                         //                                                    .writedata
		.TIMER_s1_chipselect                                       (mm_interconnect_0_timer_s1_chipselect),                        //                                                    .chipselect
		.timer_timestamp_s1_address                                (mm_interconnect_0_timer_timestamp_s1_address),                 //                                  timer_timestamp_s1.address
		.timer_timestamp_s1_write                                  (mm_interconnect_0_timer_timestamp_s1_write),                   //                                                    .write
		.timer_timestamp_s1_readdata                               (mm_interconnect_0_timer_timestamp_s1_readdata),                //                                                    .readdata
		.timer_timestamp_s1_writedata                              (mm_interconnect_0_timer_timestamp_s1_writedata),               //                                                    .writedata
		.timer_timestamp_s1_chipselect                             (mm_interconnect_0_timer_timestamp_s1_chipselect)               //                                                    .chipselect
	);

	DE0_LT24_SOPC_irq_mapper irq_mapper (
		.clk           (alt_pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),           // receiver7.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (alt_pll_c0_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (alt_pll_c0_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (alt_pll_c2_clk),                     //       receiver_clk.clk
		.sender_clk     (alt_pll_c0_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (alt_pll_c0_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver6_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (alt_pll_c0_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver7_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk            (alt_pll_c0_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (alt_pll_c2_clk),                     //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
