// MTL_SOPC.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module MTL_SOPC (
		input  wire        clk_clk,                                       //                               clk.clk
		output wire [7:0]  cyclonespi_0_spi_interface_Config,             //        cyclonespi_0_spi_interface.Config
		input  wire        cyclonespi_0_spi_interface_SPI_CS,             //                                  .SPI_CS
		input  wire        cyclonespi_0_spi_interface_SPI_SDI,            //                                  .SPI_SDI
		output wire        cyclonespi_0_spi_interface_SPI_SDO,            //                                  .SPI_SDO
		input  wire        cyclonespi_0_spi_interface_SPI_clk,            //                                  .SPI_clk
		output wire [7:0]  cyclonespi_0_spi_interface_data_out,           //                                  .data_out
		output wire        cyclonespi_0_spi_interface_data_out_enable,    //                                  .data_out_enable
		output wire        cyclonespi_0_spi_interface_spi_irq,            //                                  .spi_irq
		input  wire        from_key_export,                               //                          from_key.export
		output wire [31:0] maptransfer_map_map_line0,                     //                   maptransfer_map.map_line0
		output wire [31:0] maptransfer_map_map_line1,                     //                                  .map_line1
		output wire [31:0] maptransfer_map_map_line2,                     //                                  .map_line2
		output wire [31:0] maptransfer_map_map_line3,                     //                                  .map_line3
		output wire [31:0] maptransfer_map_map_line4,                     //                                  .map_line4
		output wire [31:0] maptransfer_map_map_line5,                     //                                  .map_line5
		output wire [31:0] maptransfer_map_map_line6,                     //                                  .map_line6
		output wire [31:0] maptransfer_map_map_line7,                     //                                  .map_line7
		input  wire [31:0] mtl_interface_irq_0_mtl_intreface_mtl_counter, // mtl_interface_irq_0_mtl_intreface.mtl_counter
		input  wire        mtl_interface_irq_0_mtl_intreface_mtl_irq,     //                                  .mtl_irq
		output wire        mtl_interface_irq_0_mtl_intreface_mtl_reset,   //                                  .mtl_reset
		output wire [3:0]  mtl_interface_irq_0_mtl_intreface_mtl_mode,    //                                  .mtl_mode
		input  wire        reset_reset_n,                                 //                             reset.reset_n
		output wire [3:0]  testled_external_connection_export,            //       testled_external_connection.export
		input  wire [19:0] touchdata_ext_export,                          //                     touchdata_ext.export
		output wire        turn_ext_export                                //                          turn_ext.export
	);

	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // CPU:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [21:0] cpu_data_master_address;                                   // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                      // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_readdatavalid;                             // mm_interconnect_0:CPU_data_master_readdatavalid -> CPU:d_readdatavalid
	wire         cpu_data_master_write;                                     // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [16:0] cpu_instruction_master_address;                            // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                               // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:CPU_instruction_master_readdatavalid -> CPU:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire   [2:0] mm_interconnect_0_maptransfer_avalon_slave_address;        // mm_interconnect_0:mapTransfer_avalon_slave_address -> mapTransfer:address
	wire         mm_interconnect_0_maptransfer_avalon_slave_write;          // mm_interconnect_0:mapTransfer_avalon_slave_write -> mapTransfer:write
	wire  [31:0] mm_interconnect_0_maptransfer_avalon_slave_writedata;      // mm_interconnect_0:mapTransfer_avalon_slave_writedata -> mapTransfer:writedata
	wire  [31:0] mm_interconnect_0_mtl_interface_irq_0_avs_s0_readdata;     // mtl_interface_irq_0:avs_s0_readdata -> mm_interconnect_0:mtl_interface_irq_0_avs_s0_readdata
	wire         mm_interconnect_0_mtl_interface_irq_0_avs_s0_waitrequest;  // mtl_interface_irq_0:avs_s0_waitrequest -> mm_interconnect_0:mtl_interface_irq_0_avs_s0_waitrequest
	wire   [7:0] mm_interconnect_0_mtl_interface_irq_0_avs_s0_address;      // mm_interconnect_0:mtl_interface_irq_0_avs_s0_address -> mtl_interface_irq_0:avs_s0_address
	wire         mm_interconnect_0_mtl_interface_irq_0_avs_s0_read;         // mm_interconnect_0:mtl_interface_irq_0_avs_s0_read -> mtl_interface_irq_0:avs_s0_read
	wire         mm_interconnect_0_mtl_interface_irq_0_avs_s0_write;        // mm_interconnect_0:mtl_interface_irq_0_avs_s0_write -> mtl_interface_irq_0:avs_s0_write
	wire  [31:0] mm_interconnect_0_mtl_interface_irq_0_avs_s0_writedata;    // mm_interconnect_0:mtl_interface_irq_0_avs_s0_writedata -> mtl_interface_irq_0:avs_s0_writedata
	wire  [31:0] mm_interconnect_0_cyclonespi_0_avs_s0_readdata;            // cycloneSPI_0:avs_s0_readdata -> mm_interconnect_0:cycloneSPI_0_avs_s0_readdata
	wire         mm_interconnect_0_cyclonespi_0_avs_s0_waitrequest;         // cycloneSPI_0:avs_s0_waitrequest -> mm_interconnect_0:cycloneSPI_0_avs_s0_waitrequest
	wire   [7:0] mm_interconnect_0_cyclonespi_0_avs_s0_address;             // mm_interconnect_0:cycloneSPI_0_avs_s0_address -> cycloneSPI_0:avs_s0_address
	wire         mm_interconnect_0_cyclonespi_0_avs_s0_read;                // mm_interconnect_0:cycloneSPI_0_avs_s0_read -> cycloneSPI_0:avs_s0_read
	wire         mm_interconnect_0_cyclonespi_0_avs_s0_write;               // mm_interconnect_0:cycloneSPI_0_avs_s0_write -> cycloneSPI_0:avs_s0_write
	wire  [31:0] mm_interconnect_0_cyclonespi_0_avs_s0_writedata;           // mm_interconnect_0:cycloneSPI_0_avs_s0_writedata -> cycloneSPI_0:avs_s0_writedata
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;          // CPU:jtag_debug_module_readdata -> mm_interconnect_0:CPU_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;       // CPU:jtag_debug_module_waitrequest -> mm_interconnect_0:CPU_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;       // mm_interconnect_0:CPU_jtag_debug_module_debugaccess -> CPU:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;           // mm_interconnect_0:CPU_jtag_debug_module_address -> CPU:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;              // mm_interconnect_0:CPU_jtag_debug_module_read -> CPU:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;        // mm_interconnect_0:CPU_jtag_debug_module_byteenable -> CPU:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;             // mm_interconnect_0:CPU_jtag_debug_module_write -> CPU:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;         // mm_interconnect_0:CPU_jtag_debug_module_writedata -> CPU:jtag_debug_module_writedata
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                         // KEY:readdata -> mm_interconnect_0:KEY_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                          // mm_interconnect_0:KEY_s1_address -> KEY:address
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:TIMER_s1_chipselect -> TIMER:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // TIMER:readdata -> mm_interconnect_0:TIMER_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:TIMER_s1_address -> TIMER:address
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:TIMER_s1_write -> TIMER:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:TIMER_s1_writedata -> TIMER:writedata
	wire         mm_interconnect_0_testled_s1_chipselect;                   // mm_interconnect_0:TESTLED_s1_chipselect -> TESTLED:chipselect
	wire  [31:0] mm_interconnect_0_testled_s1_readdata;                     // TESTLED:readdata -> mm_interconnect_0:TESTLED_s1_readdata
	wire   [1:0] mm_interconnect_0_testled_s1_address;                      // mm_interconnect_0:TESTLED_s1_address -> TESTLED:address
	wire         mm_interconnect_0_testled_s1_write;                        // mm_interconnect_0:TESTLED_s1_write -> TESTLED:write_n
	wire  [31:0] mm_interconnect_0_testled_s1_writedata;                    // mm_interconnect_0:TESTLED_s1_writedata -> TESTLED:writedata
	wire         mm_interconnect_0_mem_s1_chipselect;                       // mm_interconnect_0:mem_s1_chipselect -> mem:chipselect
	wire  [31:0] mm_interconnect_0_mem_s1_readdata;                         // mem:readdata -> mm_interconnect_0:mem_s1_readdata
	wire  [12:0] mm_interconnect_0_mem_s1_address;                          // mm_interconnect_0:mem_s1_address -> mem:address
	wire   [3:0] mm_interconnect_0_mem_s1_byteenable;                       // mm_interconnect_0:mem_s1_byteenable -> mem:byteenable
	wire         mm_interconnect_0_mem_s1_write;                            // mm_interconnect_0:mem_s1_write -> mem:write
	wire  [31:0] mm_interconnect_0_mem_s1_writedata;                        // mm_interconnect_0:mem_s1_writedata -> mem:writedata
	wire         mm_interconnect_0_mem_s1_clken;                            // mm_interconnect_0:mem_s1_clken -> mem:clken
	wire  [31:0] mm_interconnect_0_touchdata_s1_readdata;                   // TOUCHDATA:readdata -> mm_interconnect_0:TOUCHDATA_s1_readdata
	wire   [1:0] mm_interconnect_0_touchdata_s1_address;                    // mm_interconnect_0:TOUCHDATA_s1_address -> TOUCHDATA:address
<<<<<<< HEAD
	wire         mm_interconnect_0_turn_s1_chipselect;                      // mm_interconnect_0:TURN_s1_chipselect -> TURN:chipselect
	wire  [31:0] mm_interconnect_0_turn_s1_readdata;                        // TURN:readdata -> mm_interconnect_0:TURN_s1_readdata
	wire   [1:0] mm_interconnect_0_turn_s1_address;                         // mm_interconnect_0:TURN_s1_address -> TURN:address
	wire         mm_interconnect_0_turn_s1_write;                           // mm_interconnect_0:TURN_s1_write -> TURN:write_n
	wire  [31:0] mm_interconnect_0_turn_s1_writedata;                       // mm_interconnect_0:TURN_s1_writedata -> TURN:writedata
	wire         irq_mapper_receiver0_irq;                                  // mtl_interface_irq_0:ins_irq0_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // cycloneSPI_0:ins_irq0_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // JTAG_UART:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // TIMER:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_d_irq_irq;                                             // irq_mapper:sender_irq -> CPU:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [CPU:reset_n, JTAG_UART:rst_n, KEY:reset_n, TIMER:reset_n, irq_mapper:reset, mm_interconnect_0:CPU_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset]
=======
	wire         irq_mapper_receiver0_irq;                                  // mtl_interface_irq_0:ins_irq0_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // JTAG_UART:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // TIMER:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> CPU:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [CPU:reset_n, JTAG_UART:rst_n, KEY:reset_n, TIMER:reset_n, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
>>>>>>> addd119a196e0f16961ae63bce1fbb921569d96d
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [CPU:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                         // CPU:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [TESTLED:reset_n, TOUCHDATA:reset_n, TURN:reset_n, cycloneSPI_0:reset, mem:reset, mm_interconnect_0:mapTransfer_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mtl_interface_irq_0_reset_reset_bridge_in_reset_reset, mtl_interface_irq_0:reset_reset, rst_translator_001:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [mem:reset_req, rst_translator_001:reset_req_in]

	MTL_SOPC_CPU cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	MTL_SOPC_JTAG_UART jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
<<<<<<< HEAD
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
=======
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
>>>>>>> addd119a196e0f16961ae63bce1fbb921569d96d
	);

	MTL_SOPC_KEY key (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_key_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_key_s1_readdata), //                    .readdata
		.in_port  (from_key_export)                    // external_connection.export
	);

	MTL_SOPC_TESTLED testled (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_testled_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_testled_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_testled_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_testled_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_testled_s1_readdata),   //                    .readdata
		.out_port   (testled_external_connection_export)       // external_connection.export
	);

	MTL_SOPC_TIMER timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
<<<<<<< HEAD
		.irq        (irq_mapper_receiver3_irq)               //   irq.irq
=======
		.irq        (irq_mapper_receiver2_irq)               //   irq.irq
>>>>>>> addd119a196e0f16961ae63bce1fbb921569d96d
	);

	MTL_SOPC_TOUCHDATA touchdata (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_touchdata_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_touchdata_s1_readdata), //                    .readdata
		.in_port  (touchdata_ext_export)                     // external_connection.export
	);

	MTL_SOPC_TURN turn (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_turn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_turn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_turn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_turn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_turn_s1_readdata),   //                    .readdata
		.out_port   (turn_ext_export)                       // external_connection.export
	);

	MyCycloneSPI #(
		.A_Config     (8'b00000000),
		.RetreiveAddr (8'b00000001),
		.Counter      (8'b00000010),
		.PosX         (8'b00000011),
		.PosY         (8'b00000100),
		.ImagePixel_R (8'b00010010),
		.ImagePixel_G (8'b00010011),
		.ImagePixel_B (8'b00010100),
		.A_Led70      (8'b00010110)
	) cyclonespi_0 (
		.avs_s0_address     (mm_interconnect_0_cyclonespi_0_avs_s0_address),     //        avs_s0.address
		.avs_s0_read        (mm_interconnect_0_cyclonespi_0_avs_s0_read),        //              .read
		.avs_s0_readdata    (mm_interconnect_0_cyclonespi_0_avs_s0_readdata),    //              .readdata
		.avs_s0_write       (mm_interconnect_0_cyclonespi_0_avs_s0_write),       //              .write
		.avs_s0_writedata   (mm_interconnect_0_cyclonespi_0_avs_s0_writedata),   //              .writedata
		.avs_s0_waitrequest (mm_interconnect_0_cyclonespi_0_avs_s0_waitrequest), //              .waitrequest
		.clk                (clk_clk),                                           //         clock.clk
		.reset              (rst_controller_001_reset_out_reset),                //         reset.reset
		.ins_irq0_irq       (irq_mapper_receiver1_irq),                          //      ins_irq0.irq
		.Config             (cyclonespi_0_spi_interface_Config),                 // SPI_interface.Config
		.SPI_CS             (cyclonespi_0_spi_interface_SPI_CS),                 //              .SPI_CS
		.SPI_SDI            (cyclonespi_0_spi_interface_SPI_SDI),                //              .SPI_SDI
		.SPI_SDO            (cyclonespi_0_spi_interface_SPI_SDO),                //              .SPI_SDO
		.SPI_clk            (cyclonespi_0_spi_interface_SPI_clk),                //              .SPI_clk
		.data_out           (cyclonespi_0_spi_interface_data_out),               //              .data_out
		.data_out_enable    (cyclonespi_0_spi_interface_data_out_enable),        //              .data_out_enable
		.spi_irq            (cyclonespi_0_spi_interface_spi_irq)                 //              .spi_irq
	);

	mapTransfer maptransfer (
		.clock     (clk_clk),                                              //        clock.clk
		.reset     (~reset_reset_n),                                       //        reset.reset
		.map_line0 (maptransfer_map_map_line0),                            //          map.map_line0
		.map_line1 (maptransfer_map_map_line1),                            //             .map_line1
		.map_line2 (maptransfer_map_map_line2),                            //             .map_line2
		.map_line3 (maptransfer_map_map_line3),                            //             .map_line3
		.map_line4 (maptransfer_map_map_line4),                            //             .map_line4
		.map_line5 (maptransfer_map_map_line5),                            //             .map_line5
		.map_line6 (maptransfer_map_map_line6),                            //             .map_line6
		.map_line7 (maptransfer_map_map_line7),                            //             .map_line7
		.address   (mm_interconnect_0_maptransfer_avalon_slave_address),   // avalon_slave.address
		.write     (mm_interconnect_0_maptransfer_avalon_slave_write),     //             .write
		.writedata (mm_interconnect_0_maptransfer_avalon_slave_writedata)  //             .writedata
	);

	MTL_SOPC_mem mem (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_mem_s1_address),       //     s1.address
		.clken      (mm_interconnect_0_mem_s1_clken),         //       .clken
		.chipselect (mm_interconnect_0_mem_s1_chipselect),    //       .chipselect
		.write      (mm_interconnect_0_mem_s1_write),         //       .write
		.readdata   (mm_interconnect_0_mem_s1_readdata),      //       .readdata
		.writedata  (mm_interconnect_0_mem_s1_writedata),     //       .writedata
		.byteenable (mm_interconnect_0_mem_s1_byteenable),    //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)  //       .reset_req
	);

	mtl_interface_irq #(
		.mtl_reset_addr   (3'b000),
		.mtl_mode_addr    (3'b001),
		.mtl_counter_addr (3'b010)
	) mtl_interface_irq_0 (
		.avs_s0_address     (mm_interconnect_0_mtl_interface_irq_0_avs_s0_address),     //        avs_s0.address
		.avs_s0_read        (mm_interconnect_0_mtl_interface_irq_0_avs_s0_read),        //              .read
		.avs_s0_readdata    (mm_interconnect_0_mtl_interface_irq_0_avs_s0_readdata),    //              .readdata
		.avs_s0_write       (mm_interconnect_0_mtl_interface_irq_0_avs_s0_write),       //              .write
		.avs_s0_writedata   (mm_interconnect_0_mtl_interface_irq_0_avs_s0_writedata),   //              .writedata
		.avs_s0_waitrequest (mm_interconnect_0_mtl_interface_irq_0_avs_s0_waitrequest), //              .waitrequest
		.clock_clk          (clk_clk),                                                  //         clock.clk
		.reset_reset        (rst_controller_001_reset_out_reset),                       //         reset.reset
		.ins_irq0_irq       (irq_mapper_receiver0_irq),                                 //      ins_irq0.irq
<<<<<<< HEAD
		.mtl_counter        (mtl_interface_irq_0_mtl_intreface_mtl_counter),            // mtl_intreface.mtl_counter
		.mtl_irq            (mtl_interface_irq_0_mtl_intreface_mtl_irq),                //              .mtl_irq
		.mtl_reset          (mtl_interface_irq_0_mtl_intreface_mtl_reset),              //              .mtl_reset
		.mtl_mode           (mtl_interface_irq_0_mtl_intreface_mtl_mode)                //              .mtl_mode
=======
		.mtl_irq            (mtl_interface_irq_0_mtl_interface_mtl_irq),                // mtl_interface.mtl_irq
		.mtl_reset          (mtl_interface_irq_0_mtl_interface_mtl_reset),              //              .mtl_reset
		.mtl_mode           (mtl_interface_irq_0_mtl_interface_mtl_mode),               //              .mtl_mode
		.mtl_counter        (mtl_interface_irq_0_mtl_interface_mtl_counter)             //              .mtl_counter
>>>>>>> addd119a196e0f16961ae63bce1fbb921569d96d
	);

	MTL_SOPC_mm_interconnect_0 mm_interconnect_0 (
		.CLK_50_clk_clk                                        (clk_clk),                                                   //                                      CLK_50_clk.clk
		.CPU_reset_n_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                            //               CPU_reset_n_reset_bridge_in_reset.reset
		.mapTransfer_reset_reset_bridge_in_reset_reset         (rst_controller_001_reset_out_reset),                        //         mapTransfer_reset_reset_bridge_in_reset.reset
		.mtl_interface_irq_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // mtl_interface_irq_0_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address                               (cpu_data_master_address),                                   //                                 CPU_data_master.address
		.CPU_data_master_waitrequest                           (cpu_data_master_waitrequest),                               //                                                .waitrequest
		.CPU_data_master_byteenable                            (cpu_data_master_byteenable),                                //                                                .byteenable
		.CPU_data_master_read                                  (cpu_data_master_read),                                      //                                                .read
		.CPU_data_master_readdata                              (cpu_data_master_readdata),                                  //                                                .readdata
		.CPU_data_master_readdatavalid                         (cpu_data_master_readdatavalid),                             //                                                .readdatavalid
		.CPU_data_master_write                                 (cpu_data_master_write),                                     //                                                .write
		.CPU_data_master_writedata                             (cpu_data_master_writedata),                                 //                                                .writedata
		.CPU_data_master_debugaccess                           (cpu_data_master_debugaccess),                               //                                                .debugaccess
		.CPU_instruction_master_address                        (cpu_instruction_master_address),                            //                          CPU_instruction_master.address
		.CPU_instruction_master_waitrequest                    (cpu_instruction_master_waitrequest),                        //                                                .waitrequest
		.CPU_instruction_master_read                           (cpu_instruction_master_read),                               //                                                .read
		.CPU_instruction_master_readdata                       (cpu_instruction_master_readdata),                           //                                                .readdata
		.CPU_instruction_master_readdatavalid                  (cpu_instruction_master_readdatavalid),                      //                                                .readdatavalid
		.CPU_jtag_debug_module_address                         (mm_interconnect_0_cpu_jtag_debug_module_address),           //                           CPU_jtag_debug_module.address
		.CPU_jtag_debug_module_write                           (mm_interconnect_0_cpu_jtag_debug_module_write),             //                                                .write
		.CPU_jtag_debug_module_read                            (mm_interconnect_0_cpu_jtag_debug_module_read),              //                                                .read
		.CPU_jtag_debug_module_readdata                        (mm_interconnect_0_cpu_jtag_debug_module_readdata),          //                                                .readdata
		.CPU_jtag_debug_module_writedata                       (mm_interconnect_0_cpu_jtag_debug_module_writedata),         //                                                .writedata
		.CPU_jtag_debug_module_byteenable                      (mm_interconnect_0_cpu_jtag_debug_module_byteenable),        //                                                .byteenable
		.CPU_jtag_debug_module_waitrequest                     (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),       //                                                .waitrequest
		.CPU_jtag_debug_module_debugaccess                     (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),       //                                                .debugaccess
		.cycloneSPI_0_avs_s0_address                           (mm_interconnect_0_cyclonespi_0_avs_s0_address),             //                             cycloneSPI_0_avs_s0.address
		.cycloneSPI_0_avs_s0_write                             (mm_interconnect_0_cyclonespi_0_avs_s0_write),               //                                                .write
		.cycloneSPI_0_avs_s0_read                              (mm_interconnect_0_cyclonespi_0_avs_s0_read),                //                                                .read
		.cycloneSPI_0_avs_s0_readdata                          (mm_interconnect_0_cyclonespi_0_avs_s0_readdata),            //                                                .readdata
		.cycloneSPI_0_avs_s0_writedata                         (mm_interconnect_0_cyclonespi_0_avs_s0_writedata),           //                                                .writedata
		.cycloneSPI_0_avs_s0_waitrequest                       (mm_interconnect_0_cyclonespi_0_avs_s0_waitrequest),         //                                                .waitrequest
		.JTAG_UART_avalon_jtag_slave_address                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                     JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                .write
		.JTAG_UART_avalon_jtag_slave_read                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                .read
		.JTAG_UART_avalon_jtag_slave_readdata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                .readdata
		.JTAG_UART_avalon_jtag_slave_writedata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.KEY_s1_address                                        (mm_interconnect_0_key_s1_address),                          //                                          KEY_s1.address
		.KEY_s1_readdata                                       (mm_interconnect_0_key_s1_readdata),                         //                                                .readdata
		.mapTransfer_avalon_slave_address                      (mm_interconnect_0_maptransfer_avalon_slave_address),        //                        mapTransfer_avalon_slave.address
		.mapTransfer_avalon_slave_write                        (mm_interconnect_0_maptransfer_avalon_slave_write),          //                                                .write
		.mapTransfer_avalon_slave_writedata                    (mm_interconnect_0_maptransfer_avalon_slave_writedata),      //                                                .writedata
		.mem_s1_address                                        (mm_interconnect_0_mem_s1_address),                          //                                          mem_s1.address
		.mem_s1_write                                          (mm_interconnect_0_mem_s1_write),                            //                                                .write
		.mem_s1_readdata                                       (mm_interconnect_0_mem_s1_readdata),                         //                                                .readdata
		.mem_s1_writedata                                      (mm_interconnect_0_mem_s1_writedata),                        //                                                .writedata
		.mem_s1_byteenable                                     (mm_interconnect_0_mem_s1_byteenable),                       //                                                .byteenable
		.mem_s1_chipselect                                     (mm_interconnect_0_mem_s1_chipselect),                       //                                                .chipselect
		.mem_s1_clken                                          (mm_interconnect_0_mem_s1_clken),                            //                                                .clken
		.mtl_interface_irq_0_avs_s0_address                    (mm_interconnect_0_mtl_interface_irq_0_avs_s0_address),      //                      mtl_interface_irq_0_avs_s0.address
		.mtl_interface_irq_0_avs_s0_write                      (mm_interconnect_0_mtl_interface_irq_0_avs_s0_write),        //                                                .write
		.mtl_interface_irq_0_avs_s0_read                       (mm_interconnect_0_mtl_interface_irq_0_avs_s0_read),         //                                                .read
		.mtl_interface_irq_0_avs_s0_readdata                   (mm_interconnect_0_mtl_interface_irq_0_avs_s0_readdata),     //                                                .readdata
		.mtl_interface_irq_0_avs_s0_writedata                  (mm_interconnect_0_mtl_interface_irq_0_avs_s0_writedata),    //                                                .writedata
		.mtl_interface_irq_0_avs_s0_waitrequest                (mm_interconnect_0_mtl_interface_irq_0_avs_s0_waitrequest),  //                                                .waitrequest
		.TESTLED_s1_address                                    (mm_interconnect_0_testled_s1_address),                      //                                      TESTLED_s1.address
		.TESTLED_s1_write                                      (mm_interconnect_0_testled_s1_write),                        //                                                .write
		.TESTLED_s1_readdata                                   (mm_interconnect_0_testled_s1_readdata),                     //                                                .readdata
		.TESTLED_s1_writedata                                  (mm_interconnect_0_testled_s1_writedata),                    //                                                .writedata
		.TESTLED_s1_chipselect                                 (mm_interconnect_0_testled_s1_chipselect),                   //                                                .chipselect
		.TIMER_s1_address                                      (mm_interconnect_0_timer_s1_address),                        //                                        TIMER_s1.address
		.TIMER_s1_write                                        (mm_interconnect_0_timer_s1_write),                          //                                                .write
		.TIMER_s1_readdata                                     (mm_interconnect_0_timer_s1_readdata),                       //                                                .readdata
		.TIMER_s1_writedata                                    (mm_interconnect_0_timer_s1_writedata),                      //                                                .writedata
		.TIMER_s1_chipselect                                   (mm_interconnect_0_timer_s1_chipselect),                     //                                                .chipselect
		.TOUCHDATA_s1_address                                  (mm_interconnect_0_touchdata_s1_address),                    //                                    TOUCHDATA_s1.address
		.TOUCHDATA_s1_readdata                                 (mm_interconnect_0_touchdata_s1_readdata),                   //                                                .readdata
		.TURN_s1_address                                       (mm_interconnect_0_turn_s1_address),                         //                                         TURN_s1.address
		.TURN_s1_write                                         (mm_interconnect_0_turn_s1_write),                           //                                                .write
		.TURN_s1_readdata                                      (mm_interconnect_0_turn_s1_readdata),                        //                                                .readdata
		.TURN_s1_writedata                                     (mm_interconnect_0_turn_s1_writedata),                       //                                                .writedata
		.TURN_s1_chipselect                                    (mm_interconnect_0_turn_s1_chipselect)                       //                                                .chipselect
	);

	MTL_SOPC_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
<<<<<<< HEAD
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
=======
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
>>>>>>> addd119a196e0f16961ae63bce1fbb921569d96d
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
